�  �؎Ў�����f� |  ��L�� �� ��@�� �r�� ��fUf��f��f� �  f�Аf�f�                                                                                                                                                                                                                                                                                                                                                                                                                                                        U��
f� �؎Ў������م   fUf��f��gf�Eg�E�gf�E�f���g�E�gf�E�f�f�fUf��f��gf�Ugf�Eg�U�g�E�gf�U�gf�E��f�f�fUf����f]f�fUf��f��gf�Ef��g�E�gf�Eg�E�gf�Ef��g�E�gU��f�f�fUf��f�� �gf�E�gf�E�f�f�fUf��gf�E"��f]f�fUf��f��gf�Egf�E�gf�Egf�E�gf�E�gf�(�f�f�fUf��f���gf�E�����gf�Egf�Pgf�Ugf� g�E�g�}� uՐf�f�fUf��fWfVfSf��0gf�E�    fh%�  f����f��f�Ж    gf�E�    �� gf�E�gf�E�f� �  gf�]�f�   f�PAMSgf�u�f���f��gf�E�gf�M�gf�U�gf�}�PAMStfh;�  f�4���f��� gf�}�~gf�E�gf�@f��f��tSgf�E�gf�@f��u9f�Жgf�U�gf�gf�ŀ�  f�Жgf�U�gf�Rgf�ń�  f�Жf��f�Жgf�}� t��gf�E�gf�}�	�&���fhE�  f����f��gf�e�f[f^f_f]f�fUf��f��f�����fh�   f����f��g�E�gf�E�f��f��fPfh�   f����f��f�`�  fjfPf����f��f�����gf�E�gf�E�f��fPf�����f��f��  fPfjf�����f���f�f�fUf��fhK�  f�����f��f����f�M�����U����Ef�E��E���E��E���U����Ef�E��E��f�f�E��E���U����U�Ef�U��E��U��E����U��S��h�   h�  ��������E����Ph�  �������E����Ph�  ������j h�  ������j h�  �������E��Ph�  �k������E��Ph�  �W������E����Ph�  �@������E����Ph�  �)�����j$h�  �������E�E��J�h�  ���������%�   ��u��E�    ��]��C�E�h�  ������f��E��}��   ~ڋE�P��U�����]���U��� �E�E�E�� <u!�E��@<Eu�E��@<Lu�E��@<Ft
�    ��   �E�    �   �E�P�EE���ЉE�E� ����   �E�P�EЉE��E�@�E��E�    ��U��B�E��E�H�M����E��E�P�E�9�w؋E�P�E�@ЉE��E�    ��E�P�U��  �E��E�P�E�@)E�9�w����E��E��@,��9E��;����E�@��U����U���h   h�  jd������h   �������E�}� u
j���������E��h��  �Ѓ���try to detect memory: failed.
 ok.
 ....loading.....
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ��   �� ��   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ELF                 4   �      4    (               i  �8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �t$��
  �   f� �؎Ў����輐8 ��
  j j�`��T�\  ����a���j j `��T�S  ����a���j j`��T�J  ����a���j j`��T�A  ����a���j j`��T�8  ����a���j j`��T�/  ����a���j j`��T�&  ����a���j j`��T�  ����a���j j`��T�  ����a���j`��T�  ����a���j
`��T�  ����a���j`��T��  ����a���j`��T��  ����a���j`��T��  ����a���j`��T��  ����a���j j`��T��  ����a���j`��T��  ����a���j j`��T��  ����a���j j`��T��  ����a���j j`��T�  ����a���j j `��T�  ����a���U����E��f�E��Ef�E��E��f�E�U����U����Ef�E�E����� �E��}�� vf�M� ��E���E�E�E�f��E�E�f�P�E���E��P�E����f% fE�E�f�P�E���E��P���U����U�Ef�U�f�E��E�Ef��E�U�f�P�E�U�f�P�E���Ef�P���U����E�    ��E���j j j P�������E��}��   ~�h��  j�j j�������h��  j�j j��������� h   P���������U�������]�U����Ef�E��E���E��E���U����U�Ef�U��E��U��E����U����]�U����]�U����E��f�E��Ef�E��E��f�E�]����U����]�U���������U��h�
 �u����������U��h �u����������U��h �u���������U��h- �u���������U��h< �u���������U��hH �u�x��������U��hR �u�b��������U��hh �u�L��������U��hx �u�6��������U��h� �u� ��������U��h� �u�
��������U��h� �u����������U��h� �u����������U��h� �u����������U��h� �u���������U��h� �u���������U��h �u���������U��h! �u�p��������U��h0 �u�Z��������U��hO �u�D��������U��jj �������j j!�������jj!������jj!������jh�   ������j(h�   ������jh�   ������jh�   �v�����h�   j!�g�����h�   h�   �U��������U��m �}~j h�   �6�����j j �*��������U����E�    �%�(  �E���� h �  RjP�������E��}�vՃ�hG  j �e  ����hf  j�S  ����h�  j�A  ����h�  j�/  ����h�  j�  ����h�  j�  ����h j��   ����h  j��   ����h? j��   ����h\ j
��   ����hy j�   ����h� j�   ����h� j�   ����h� j�{   ����h� j�i   ����h j�W   ����h) j�E   ����hH j�3   ����hg j�!   ���� ��h   P�������������U����}~������%�E�U��� h �  PjR�j������    ��U��S���}~x�m �}2j!�������E�   �������!ЈE��E�Pj!��������=�mh�   ��������E�   �������!ЈE��E�Ph�   ���������]���U��S���}~t�m �}0j!�v������ËE�   �����	؈E��E�Pj!�o������;�mh�   �?������ËE�   �����	؈E��E�Ph�   �5��������]���U���A����]�U���=����]�U����U�Ef�U��E��U��E����U����� ���� ��j ���������U����E��.  j6jC�������E���Pj@�������E�����Pj@��������h� j ��������j �<��������U�����     �������U����E�� ����������������U����  Unknown exception. Device Error. Debug Exception NMI Interrupt. Breakpoint. Overflow. BOUND Range Exceeded. Invalid Opcode. Device Not Available. Double Fault. Invalid TSS Segment Not Present. Stack-Segment Fault. General Protection. Page Fault. X87 FPU Floating Point Error. Alignment Check. Machine Check. SIMD Floating Point Exception. Virtualization Exception. GCC: (GNU) 7.1.0  .shstrtab .text .rodata .bss .comment                                                           �
                          �
 �  m                          � i  ,                        0       i                                 z  '                  